-- my_nios1_slave_template_1.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity my_nios1_slave_template_1 is
	generic (
		DATA_WIDTH          : integer := 32;
		ENABLE_SYNC_SIGNALS : integer := 0;
		MODE_0              : integer := 1;
		MODE_1              : integer := 1;
		MODE_2              : integer := 1;
		MODE_3              : integer := 1;
		MODE_4              : integer := 1;
		MODE_5              : integer := 1;
		MODE_6              : integer := 1;
		MODE_7              : integer := 1;
		MODE_8              : integer := 1;
		MODE_9              : integer := 1;
		MODE_10             : integer := 1;
		MODE_11             : integer := 1;
		MODE_12             : integer := 1;
		MODE_13             : integer := 1;
		MODE_14             : integer := 1;
		MODE_15             : integer := 1;
		IRQ_EN              : integer := 0
	);
	port (
		clk              : in  std_logic                     := '0';             --       clock_reset.clk
		reset            : in  std_logic                     := '0';             -- clock_reset_reset.reset
		slave_address    : in  std_logic_vector(8 downto 0)  := (others => '0'); --                s0.address
		slave_read       : in  std_logic                     := '0';             --                  .read
		slave_write      : in  std_logic                     := '0';             --                  .write
		slave_readdata   : out std_logic_vector(31 downto 0);                    --                  .readdata
		slave_writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => '0'); --                  .byteenable
		user_datain_0    : in  std_logic_vector(31 downto 0) := (others => '0'); --    user_interface.export
		user_datain_1    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_2    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_3    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_4    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_5    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_6    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_7    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_8    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_9    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_10   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_11   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_12   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_13   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_14   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		user_datain_15   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .export
		slave_irq        : out std_logic;
		user_chipselect  : out std_logic_vector(15 downto 0);
		user_dataout_0   : out std_logic_vector(31 downto 0);
		user_dataout_1   : out std_logic_vector(31 downto 0);
		user_dataout_10  : out std_logic_vector(31 downto 0);
		user_dataout_11  : out std_logic_vector(31 downto 0);
		user_dataout_12  : out std_logic_vector(31 downto 0);
		user_dataout_13  : out std_logic_vector(31 downto 0);
		user_dataout_14  : out std_logic_vector(31 downto 0);
		user_dataout_15  : out std_logic_vector(31 downto 0);
		user_dataout_2   : out std_logic_vector(31 downto 0);
		user_dataout_3   : out std_logic_vector(31 downto 0);
		user_dataout_4   : out std_logic_vector(31 downto 0);
		user_dataout_5   : out std_logic_vector(31 downto 0);
		user_dataout_6   : out std_logic_vector(31 downto 0);
		user_dataout_7   : out std_logic_vector(31 downto 0);
		user_dataout_8   : out std_logic_vector(31 downto 0);
		user_dataout_9   : out std_logic_vector(31 downto 0);
		user_read        : out std_logic;
		user_write       : out std_logic
	);
end entity my_nios1_slave_template_1;

architecture rtl of my_nios1_slave_template_1 is
	component slave_template is
		generic (
			DATA_WIDTH          : integer := 32;
			ENABLE_SYNC_SIGNALS : integer := 0;
			MODE_0              : integer := 2;
			MODE_1              : integer := 2;
			MODE_2              : integer := 2;
			MODE_3              : integer := 2;
			MODE_4              : integer := 2;
			MODE_5              : integer := 2;
			MODE_6              : integer := 2;
			MODE_7              : integer := 2;
			MODE_8              : integer := 2;
			MODE_9              : integer := 2;
			MODE_10             : integer := 2;
			MODE_11             : integer := 2;
			MODE_12             : integer := 2;
			MODE_13             : integer := 2;
			MODE_14             : integer := 2;
			MODE_15             : integer := 2;
			IRQ_EN              : integer := 0
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			slave_address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			slave_read       : in  std_logic                     := 'X';             -- read
			slave_write      : in  std_logic                     := 'X';             -- write
			slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			slave_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			user_datain_0    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_1    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_2    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_3    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_4    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_5    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_6    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_7    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_8    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_9    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_10   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_11   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_12   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_13   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_14   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_15   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			slave_irq        : out std_logic;                                        -- irq
			user_dataout_0   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_1   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_2   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_3   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_4   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_5   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_6   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_7   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_8   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_9   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_10  : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_11  : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_12  : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_13  : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_14  : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_15  : out std_logic_vector(31 downto 0);                    -- export
			user_write       : out std_logic;                                        -- export
			user_read        : out std_logic;                                        -- export
			user_chipselect  : out std_logic_vector(15 downto 0)                     -- export
		);
	end component slave_template;

begin

	slave_template_1 : component slave_template
		generic map (
			DATA_WIDTH          => DATA_WIDTH,
			ENABLE_SYNC_SIGNALS => ENABLE_SYNC_SIGNALS,
			MODE_0              => MODE_0,
			MODE_1              => MODE_1,
			MODE_2              => MODE_2,
			MODE_3              => MODE_3,
			MODE_4              => MODE_4,
			MODE_5              => MODE_5,
			MODE_6              => MODE_6,
			MODE_7              => MODE_7,
			MODE_8              => MODE_8,
			MODE_9              => MODE_9,
			MODE_10             => MODE_10,
			MODE_11             => MODE_11,
			MODE_12             => MODE_12,
			MODE_13             => MODE_13,
			MODE_14             => MODE_14,
			MODE_15             => MODE_15,
			IRQ_EN              => IRQ_EN
		)
		port map (
			clk              => clk,              --       clock_reset.clk
			reset            => reset,            -- clock_reset_reset.reset
			slave_address    => slave_address,    --                s0.address
			slave_read       => slave_read,       --                  .read
			slave_write      => slave_write,      --                  .write
			slave_readdata   => slave_readdata,   --                  .readdata
			slave_writedata  => slave_writedata,  --                  .writedata
			slave_byteenable => slave_byteenable, --                  .byteenable
			user_datain_0    => user_datain_0,    --    user_interface.export
			user_datain_1    => user_datain_1,    --                  .export
			user_datain_2    => user_datain_2,    --                  .export
			user_datain_3    => user_datain_3,    --                  .export
			user_datain_4    => user_datain_4,    --                  .export
			user_datain_5    => user_datain_5,    --                  .export
			user_datain_6    => user_datain_6,    --                  .export
			user_datain_7    => user_datain_7,    --                  .export
			user_datain_8    => user_datain_8,    --                  .export
			user_datain_9    => user_datain_9,    --                  .export
			user_datain_10   => user_datain_10,   --                  .export
			user_datain_11   => user_datain_11,   --                  .export
			user_datain_12   => user_datain_12,   --                  .export
			user_datain_13   => user_datain_13,   --                  .export
			user_datain_14   => user_datain_14,   --                  .export
			user_datain_15   => user_datain_15,   --                  .export
			slave_irq        => open,             --       (terminated)
			user_dataout_0   => open,             --       (terminated)
			user_dataout_1   => open,             --       (terminated)
			user_dataout_2   => open,             --       (terminated)
			user_dataout_3   => open,             --       (terminated)
			user_dataout_4   => open,             --       (terminated)
			user_dataout_5   => open,             --       (terminated)
			user_dataout_6   => open,             --       (terminated)
			user_dataout_7   => open,             --       (terminated)
			user_dataout_8   => open,             --       (terminated)
			user_dataout_9   => open,             --       (terminated)
			user_dataout_10  => open,             --       (terminated)
			user_dataout_11  => open,             --       (terminated)
			user_dataout_12  => open,             --       (terminated)
			user_dataout_13  => open,             --       (terminated)
			user_dataout_14  => open,             --       (terminated)
			user_dataout_15  => open,             --       (terminated)
			user_write       => open,             --       (terminated)
			user_read        => open,             --       (terminated)
			user_chipselect  => open              --       (terminated)
		);

end architecture rtl; -- of my_nios1_slave_template_1
